//created by Joonseo Park

`ifndef AUDIO_PARAMS
`define AUDIO_PARAMS

//parameter START_ADDR = 32'h0000AF30;
//parameter END_ADDR = 32'h000700A0;

//parameter START_ADDR = 0;
//parameter END_ADDR = 32'h0000B780;

`endif